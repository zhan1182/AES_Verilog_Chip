library verilog;
use verilog.vl_types.all;
entity tb_inv_mix_column is
end tb_inv_mix_column;
